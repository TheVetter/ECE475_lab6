-- Name 
-- Student ID 

-- TODO: Do all of lab

